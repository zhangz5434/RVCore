Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;

Entity Decoder5_32 is
	Port(
		SELECTOR : IN std_logic_vector(4 downto 0);
		SELECTED : OUT std_logic_vector(31 downto 0)
	);
End Entity Decoder5_32;

Architecture Behavioral of Decoder5_32 is 
Begin
	Process(SELECTOR) is
	Begin
		case SELECTOR is
			when "00000" =>
				SELECTED <= "00000000000000000000000000000001";
			when "00001" =>
				SELECTED <= "00000000000000000000000000000010";
			when "00010" =>
				SELECTED <= "00000000000000000000000000000100";
			when "00011" =>
				SELECTED <= "00000000000000000000000000001000";
			when "00100" =>
				SELECTED <= "00000000000000000000000000010000";
			when "00101" =>
				SELECTED <= "00000000000000000000000000100000";
			when "00110" =>
				SELECTED <= "00000000000000000000000001000000";
			when "00111" =>
				SELECTED <= "00000000000000000000000010000000";
			when "01000" =>
				SELECTED <= "00000000000000000000000100000000";
			when "01001" =>
				SELECTED <= "00000000000000000000001000000000";
			when "01010" =>
				SELECTED <= "00000000000000000000010000000000";
			when "01011" =>
				SELECTED <= "00000000000000000000100000000000";
			when "01100" =>
				SELECTED <= "00000000000000000001000000000000";
			when "01101" =>
				SELECTED <= "00000000000000000010000000000000";
			when "01110" =>
				SELECTED <= "00000000000000000100000000000000";
			when "01111" =>
				SELECTED <= "00000000000000001000000000000000";
			when "10000" =>
				SELECTED <= "00000000000000010000000000000000";
			when "10001" =>
				SELECTED <= "00000000000000100000000000000000";
			when "10010" =>
				SELECTED <= "00000000000001000000000000000000";
			when "10011" =>
				SELECTED <= "00000000000010000000000000000000";
			when "10100" =>
				SELECTED <= "00000000000100000000000000000000";
			when "10101" =>
				SELECTED <= "00000000001000000000000000000000";
			when "10110" =>
				SELECTED <= "00000000010000000000000000000000";
			when "10111" =>
				SELECTED <= "00000000100000000000000000000000";
			when "11000" =>
				SELECTED <= "00000001000000000000000000000000";
			when "11001" =>
				SELECTED <= "00000010000000000000000000000000";
			when "11010" =>
				SELECTED <= "00000100000000000000000000000000";
			when "11011" =>
				SELECTED <= "00001000000000000000000000000000";
			when "11100" =>
				SELECTED <= "00010000000000000000000000000000";
			when "11101" =>
				SELECTED <= "00100000000000000000000000000000";
			when "11110" =>
				SELECTED <= "01000000000000000000000000000000";
			when "11111" =>
				SELECTED <= "10000000000000000000000000000000";
			when others =>
				SELECTED <= "00000000000000000000000000000000";
		end case;
	End Process;
	
End Architecture Behavioral;